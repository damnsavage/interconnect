module bin_mux_casez(valids_r, current_idx);
   input [`NUM_SINKS-1:0] valids_r; 

   output [`LOG2_NUM_SINKS-1:0] current_idx;
   reg    [`LOG2_NUM_SINKS-1:0] current_idx;

   always @(valids_r)
   begin
      // Needs to be manually updated when NUM_SINKS changes!!!!    
      casez (valids_r)
          // Unfortunately '?' does not work in hex
          64'b???????????????????????????????????????????????????????????????1 : current_idx = 0;
          64'b??????????????????????????????????????????????????????????????10 : current_idx = 1;
          64'b?????????????????????????????????????????????????????????????100 : current_idx = 2;
          64'b????????????????????????????????????????????????????????????1000 : current_idx = 3;
          64'b???????????????????????????????????????????????????????????10000 : current_idx = 4;
          64'b??????????????????????????????????????????????????????????100000 : current_idx = 5;
          64'b?????????????????????????????????????????????????????????1000000 : current_idx = 6;
          64'b????????????????????????????????????????????????????????10000000 : current_idx = 7;
          64'b???????????????????????????????????????????????????????100000000 : current_idx = 8;
          64'b??????????????????????????????????????????????????????1000000000 : current_idx = 9;
          64'b?????????????????????????????????????????????????????10000000000 : current_idx = 10;
          64'b????????????????????????????????????????????????????100000000000 : current_idx = 11;
          64'b???????????????????????????????????????????????????1000000000000 : current_idx = 12;
          64'b??????????????????????????????????????????????????10000000000000 : current_idx = 13;
          64'b?????????????????????????????????????????????????100000000000000 : current_idx = 14;
          64'b????????????????????????????????????????????????1000000000000000 : current_idx = 15;
          64'b???????????????????????????????????????????????10000000000000000 : current_idx = 16;
          64'b??????????????????????????????????????????????100000000000000000 : current_idx = 17;
          64'b?????????????????????????????????????????????1000000000000000000 : current_idx = 18;
          64'b????????????????????????????????????????????10000000000000000000 : current_idx = 19;
          64'b???????????????????????????????????????????100000000000000000000 : current_idx = 20;
          64'b??????????????????????????????????????????1000000000000000000000 : current_idx = 21;
          64'b?????????????????????????????????????????10000000000000000000000 : current_idx = 22;
          64'b????????????????????????????????????????100000000000000000000000 : current_idx = 23;
          64'b???????????????????????????????????????1000000000000000000000000 : current_idx = 24;
          64'b??????????????????????????????????????10000000000000000000000000 : current_idx = 25;
          64'b?????????????????????????????????????100000000000000000000000000 : current_idx = 26;
          64'b????????????????????????????????????1000000000000000000000000000 : current_idx = 27;
          64'b???????????????????????????????????10000000000000000000000000000 : current_idx = 28;
          64'b??????????????????????????????????100000000000000000000000000000 : current_idx = 29;
          64'b?????????????????????????????????1000000000000000000000000000000 : current_idx = 30;
          64'b????????????????????????????????10000000000000000000000000000000 : current_idx = 31;
          64'b???????????????????????????????100000000000000000000000000000000 : current_idx = 32;
          64'b??????????????????????????????1000000000000000000000000000000000 : current_idx = 33;
          64'b?????????????????????????????10000000000000000000000000000000000 : current_idx = 34;
          64'b????????????????????????????100000000000000000000000000000000000 : current_idx = 35;
          64'b???????????????????????????1000000000000000000000000000000000000 : current_idx = 36;
          64'b??????????????????????????10000000000000000000000000000000000000 : current_idx = 37;
          64'b?????????????????????????100000000000000000000000000000000000000 : current_idx = 38;
          64'b????????????????????????1000000000000000000000000000000000000000 : current_idx = 39;
          64'b???????????????????????10000000000000000000000000000000000000000 : current_idx = 40;
          64'b??????????????????????100000000000000000000000000000000000000000 : current_idx = 41;
          64'b?????????????????????1000000000000000000000000000000000000000000 : current_idx = 42;
          64'b????????????????????10000000000000000000000000000000000000000000 : current_idx = 43;
          64'b???????????????????100000000000000000000000000000000000000000000 : current_idx = 44;
          64'b??????????????????1000000000000000000000000000000000000000000000 : current_idx = 45;
          64'b?????????????????10000000000000000000000000000000000000000000000 : current_idx = 46;
          64'b????????????????100000000000000000000000000000000000000000000000 : current_idx = 47;
          64'b???????????????1000000000000000000000000000000000000000000000000 : current_idx = 48;
          64'b??????????????10000000000000000000000000000000000000000000000000 : current_idx = 49;
          64'b?????????????100000000000000000000000000000000000000000000000000 : current_idx = 50;
          64'b????????????1000000000000000000000000000000000000000000000000000 : current_idx = 51;
          64'b???????????10000000000000000000000000000000000000000000000000000 : current_idx = 52;
          64'b??????????100000000000000000000000000000000000000000000000000000 : current_idx = 53;
          64'b?????????1000000000000000000000000000000000000000000000000000000 : current_idx = 54;
          64'b????????10000000000000000000000000000000000000000000000000000000 : current_idx = 55;
          64'b???????100000000000000000000000000000000000000000000000000000000 : current_idx = 56;
          64'b??????1000000000000000000000000000000000000000000000000000000000 : current_idx = 57;
          64'b?????10000000000000000000000000000000000000000000000000000000000 : current_idx = 58;
          64'b????100000000000000000000000000000000000000000000000000000000000 : current_idx = 59;
          64'b???1000000000000000000000000000000000000000000000000000000000000 : current_idx = 60;
          64'b??10000000000000000000000000000000000000000000000000000000000000 : current_idx = 61;
          64'b?100000000000000000000000000000000000000000000000000000000000000 : current_idx = 62;
          64'b1000000000000000000000000000000000000000000000000000000000000000 : current_idx = 63;
//          64'h???????????????1 : current_idx = 0;
//          64'h???????????????2 : current_idx = 1;
//          64'h???????????????4 : current_idx = 2;
//          64'h???????????????8 : current_idx = 3;
//          64'h??????????????10 : current_idx = 4;
//          64'h??????????????20 : current_idx = 5;
//          64'h??????????????40 : current_idx = 6;
//          64'h??????????????80 : current_idx = 7;
//          64'h?????????????100 : current_idx = 8;
//          64'h?????????????200 : current_idx = 9;
//          64'h?????????????400 : current_idx = 10;
//          64'h?????????????800 : current_idx = 11;
//          64'h????????????1000 : current_idx = 12;
//          64'h????????????2000 : current_idx = 13;
//          64'h????????????4000 : current_idx = 14;
//          64'h????????????8000 : current_idx = 15;
//          64'h???????????10000 : current_idx = 16;
//          64'h???????????20000 : current_idx = 17;
//          64'h???????????40000 : current_idx = 18;
//          64'h???????????80000 : current_idx = 19;
//          64'h??????????100000 : current_idx = 20;
//          64'h??????????200000 : current_idx = 21;
//          64'h??????????400000 : current_idx = 22;
//          64'h??????????800000 : current_idx = 23;
//          64'h?????????1000000 : current_idx = 24;
//          64'h?????????2000000 : current_idx = 25;
//          64'h?????????4000000 : current_idx = 26;
//          64'h?????????8000000 : current_idx = 27;
//          64'h????????10000000 : current_idx = 28;
//          64'h????????20000000 : current_idx = 29;
//          64'h????????40000000 : current_idx = 30;
//          64'h????????80000000 : current_idx = 31;
//          64'h???????100000000 : current_idx = 32;
//          64'h???????200000000 : current_idx = 33;
//          64'h???????400000000 : current_idx = 34;
//          64'h???????800000000 : current_idx = 35;
//          64'h??????1000000000 : current_idx = 36;
//          64'h??????2000000000 : current_idx = 37;
//          64'h??????4000000000 : current_idx = 38;
//          64'h??????8000000000 : current_idx = 39;
//          64'h?????10000000000 : current_idx = 40;
//          64'h?????20000000000 : current_idx = 41;
//          64'h?????40000000000 : current_idx = 42;
//          64'h?????80000000000 : current_idx = 43;
//          64'h????100000000000 : current_idx = 44;
//          64'h????200000000000 : current_idx = 45;
//          64'h????400000000000 : current_idx = 46;
//          64'h????800000000000 : current_idx = 47;
//          64'h???1000000000000 : current_idx = 48;
//          64'h???2000000000000 : current_idx = 49;
//          64'h???4000000000000 : current_idx = 50;
//          64'h???8000000000000 : current_idx = 51;
//          64'h??10000000000000 : current_idx = 52;
//          64'h??20000000000000 : current_idx = 53;
//          64'h??40000000000000 : current_idx = 54;
//          64'h??80000000000000 : current_idx = 55;
//          64'h?100000000000000 : current_idx = 56;
//          64'h?200000000000000 : current_idx = 57;
//          64'h?400000000000000 : current_idx = 58;
//          64'h?800000000000000 : current_idx = 59;
//          64'h1000000000000000 : current_idx = 60;
//          64'h2000000000000000 : current_idx = 61;
//          64'h4000000000000000 : current_idx = 62;
//          64'h8000000000000000 : current_idx = 63;
          default : current_idx = 0;
      endcase
   end

endmodule



// Synthesis Results:
// synthesize -effort low -to_mapped
//
// Incremental optimization status
// ===============================
//                                     Worst - - DRC Totals - -
//                            Total  Weighted    Max       Max
// Operation                   Area  Neg Slk    Trans      Cap
// -------------------------------------------------------------------------------
//  init_iopt                  1707        0         0        0
// 
// Incremental optimization status
// ===============================
//                                     Worst - - DRC Totals - -
//                            Total  Weighted    Max       Max
// Operation                   Area  Neg Slk    Trans      Cap
// -------------------------------------------------------------------------------
//  init_delay                 1707        0         0        0
//
// delay 433 ps
//
//     Instance      Cells  Cell Area  Net Area  Total Area  Wireload
// -----------------------------------------------------------------------
// bin_mux_casez    148       1707         0        1707    <none> (D)
// 
//   Type   Instances   Area   Area %
// -----------------------------------
// inverter        29  152.044    8.9
// logic          119 1554.513   91.1
// -----------------------------------
// total          148 1706.556  100.0

// with synthesis effort high
//   Type   Instances   Area   Area %
// -----------------------------------
// inverter        20  104.858    7.8
// logic          103 1239.940   92.2
// -----------------------------------
// total          123 1344.798  100.0
